module Adc(
    input i_rst,
    input i_clk,
    output [7:0] o_data,

    output wire o_adc_clk,
    input wire [7:0] i_adc_data
);



endmodule